LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
 
LIBRARY WORK;
USE WORK.ALL;

ENTITY TB_UART_TX IS
END ENTITY;

ARCHITECTURE TEST OF TB_UART_TX IS

	COMPONENT UART_TX IS
	PORT(	DATA: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			SEND: IN STD_LOGIC;
			CLK: IN STD_LOGIC;
			ARST: IN STD_LOGIC;
			R232_TX: OUT STD_LOGIC;
			IDLE: OUT STD_LOGIC);
	END COMPONENT;
	
	SIGNAL DATA: STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL SEND: STD_LOGIC;
	SIGNAL CLK: STD_LOGIC:='0';
	SIGNAL ARST: STD_LOGIC;
	SIGNAL R232_TX: STD_LOGIC;
	SIGNAL IDLE: STD_LOGIC;
	
	CONSTANT PERIOD: TIME:= 10 NS;
	
BEGIN

	DUT: UART_TX PORT MAP(DATA, SEND, CLK, ARST, R232_TX, IDLE);
	CLK <= NOT CLK AFTER PERIOD;
	
	PROCESS IS
	BEGIN
		
		ARST <= '0';
		DATA <= "01010101";
		WAIT FOR 100 NS;
		SEND <= '1';
		WAIT FOR 200 NS;
		SEND <= '0';
		WAIT FOR 3000000 NS;
		
		DATA <= "10010001";
		wait for 100 ns;
		SEND <= '1';
		WAIT FOR 200 NS;
		SEND <= '0';
		WAIT FOR 3000000 NS;
		
	END PROCESS;
	
END TEST;